import uvm_pkg::*;
`include "uvm_macros.svh"
`include "./input_if.sv"
`include "./output_if.sv"
`include "./tr_in.sv"
`include "./tr_out.sv"
`include "./sequence_in.sv"
`include "./driver_in.sv"
`include "./driver_out.sv"
`include "./monitor_in.sv"
`include "./monitor_out.sv"
`include "./agent_in.sv"
`include "./agent_out.sv"
`include "./refmod.sv"
`include "./scoreboard.sv"
`include "./env.sv"
`include "./simple_test.sv"
